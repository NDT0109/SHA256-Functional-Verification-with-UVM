class msg_seq_item extends uvm_sequence_item;
   `uvm_object_utils(msg_seq_item)
  bit [511:0] message_single = 512'h61626380000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018; 
  bit [511:0] message_double_first = 512'h6162636462636465636465666465666765666768666768696768696A68696A6B696A6B6C6A6B6C6D6B6C6D6E6C6D6E6F6D6E6F706E6F70718000000000000000;
  bit [511:0] message_double_last = 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001C0;
  bit [511:0] messagetmp = 512'h0;
  bit msg_valid;
  bit msg_nxt;
  bit [255:0] hash;
  
   function new(string name = "msg_seq_item");
      super.new(name);
   endfunction 
endclass 
