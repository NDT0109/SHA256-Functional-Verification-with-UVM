class sha_subs extends uvm_subscriber #(msg_seq_item);


  	msg_seq_item req;
  
	`uvm_component_utils(sha_subs)
  
	
 	
	
	covergroup cg;

      	option.per_instance = 1;		
      
		BLOCK : coverpoint req.message; /*{
		option.weight = 0;
		bins message_bins[]={
	512'h2f51512a0e3108017d0b440d143a3d4a433f3d665f673b3a644d3b53102d057c6d6a684a2b074e5b30132c1e057f800000000000000000000000000000000170,
512'h34295653707916800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000038,
512'h79595b4d0c1c607f6f4f3907735f6b16247f08487f2800506e277c0945487f446e4f7408281e4a0d307347061580000000000000000000000000000000000168,
512'h58776d7429574e3860746f4269700a39374e7c3262332815281f742f8000000000000000000000000000000000000000000000000000000000000000000000e0,
512'h2961661360340f32761c247f3c5162333d42577d80000000000000000000000000000000000000000000000000000000000000000000000000000000000000a0,
512'h6c6102524d77197863456c055510334b10536e1219331768038000000000000000000000000000000000000000000000000000000000000000000000000000c8,
512'h5a508000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010,
512'h0b221e3567611841556f176f44671d7c2b49366a17051230474d206e770f443528052e8000000000000000000000000000000000000000000000000000000118,
512'h7701722d564b08552e80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000048,
512'h5860713b44654005243c725e7e3b4d426a77046880000000000000000000000000000000000000000000000000000000000000000000000000000000000000a0
};
}*/
		/*Init : coverpoint req.msg_valid; {
		option.weight = 0;
		bins msg_valid_bins[]={1
};
}*/
		/*Next : coverpoint req.msg_nxt; {
		option.weight = 0;
		bins msg_nxt_bins[]={0
};
}*/
		Digest : coverpoint req.hash; 	
	endgroup: cg
  
  
  
  	 function new(input string name = "sha_subs", uvm_component parent = null); 
		super.new(name, parent);
        req = msg_seq_item::type_id::create("req");
        cg = new();		
  	endfunction: new
  





	virtual function void write(input msg_seq_item t);

		`uvm_info(get_type_name(),"Data rcvd from Monitor ap", UVM_NONE)
		t.print();							// just print transctions

      	req = t;							// data container req
		
      cg.sample();							// sample coverage whenever received an objects from ap

		`uvm_info(get_type_name(), $sformatf(" ---- Coverage is %0f", cg.get_coverage()), UVM_NONE)  // %f -> real number in decimal format

		
	endfunction : write

	


endclass          
